/*
	Top level test module
	Instantiate every sub-test module
*/
module testCpu;
	test4Core_xori				test0();  // Test XORI on four cores
	test4Core_Addition 			test1();  // Test ADD on four cores
	test4Core_jump				test2();  // Test J on four cores
	test4Core_Subtraction 		test3();  // Test SUB on four cores
	test4Core_LoadWord			test4();  // Test LW on four cores
	test4Core_StoreWord			test5();  // Test SW on four cores
	test4Core_JumpRegister		test6();  // Test JR on four cores
	test4Core_JumpAndLink		test7();  // Test JAL on four cores
	test4Core_BranchNotEqual	test8();  // Test BNE on four cores
	test4Core_SignedLessThan	test9();  // Test SLT on four cores
	test4Core_BranchEqual		test10(); // Test BEQ on four cores
endmodule